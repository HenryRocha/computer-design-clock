LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;

ENTITY memoriaROM IS
    GENERIC (
        dataWidth : NATURAL := 8;
        addrWidth : NATURAL := 3
    );
    PORT (
        Endereco : IN std_logic_vector (addrWidth - 1 DOWNTO 0);
        Dado     : OUT std_logic_vector (dataWidth - 1 DOWNTO 0)
    );
END ENTITY;

ARCHITECTURE assincrona OF memoriaROM IS
    TYPE blocoMemoria IS ARRAY(0 TO 2 ** addrWidth - 1) OF std_logic_vector(dataWidth - 1 DOWNTO 0);

    FUNCTION initMemory
        RETURN blocoMemoria IS VARIABLE tmp : blocoMemoria := (OTHERS => (OTHERS => '0'));
    BEGIN
        tmp(0)  := "0110" & "000" & "000000000000";
        tmp(1)  := "0110" & "001" & "000000000000";
        tmp(2)  := "0110" & "010" & "000000000000";
        tmp(3)  := "0101" & "000" & "100000000000";
        tmp(4)  := "0101" & "001" & "100000000001";
        tmp(5)  := "0101" & "010" & "100000000010";
        tmp(6)  := "0100" & "111" & "010000000001";
        tmp(7)  := "0101" & "000" & "100000000000";
        tmp(8)  := "0101" & "001" & "100000000001";
        tmp(9)  := "0101" & "010" & "100000000010";
        tmp(10) := "0100" & "111" & "010000000000";
        tmp(11) := "0111" & "111" & "000000000001";
        tmp(12) := "1000" & "000" & "000000001110";
        tmp(13) := "1010" & "000" & "000000000111";
        tmp(14) := "0100" & "111" & "010000000001";
        tmp(15) := "0100" & "100" & "000000000001";
        tmp(16) := "0111" & "100" & "000000000001";
        tmp(17) := "1000" & "000" & "000000100111";
        tmp(18) := "0001" & "000" & "000000000001";
        tmp(19) := "0111" & "000" & "000000111100";
        tmp(20) := "1000" & "000" & "000000010110";
        tmp(21) := "1010" & "000" & "000000000111";
        tmp(22) := "0110" & "000" & "000000000000";
        tmp(23) := "0001" & "001" & "000000000001";
        tmp(24) := "0111" & "001" & "000000111100";
        tmp(25) := "1000" & "000" & "000000011011";
        tmp(26) := "1010" & "000" & "000000000111";
        tmp(27) := "0110" & "001" & "000000000000";
        tmp(28) := "0001" & "010" & "000000000001";
        tmp(29) := "0111" & "010" & "000000011000";
        tmp(30) := "1000" & "000" & "000000100000";
        tmp(31) := "1010" & "000" & "000000000111";
        tmp(32) := "0110" & "000" & "000000000000";
        tmp(33) := "0110" & "001" & "000000000000";
        tmp(34) := "0110" & "010" & "000000000000";
        tmp(35) := "0101" & "000" & "100000000000";
        tmp(36) := "0101" & "001" & "100000000001";
        tmp(37) := "0101" & "010" & "100000000010";
        tmp(38) := "1010" & "000" & "000000000111";
        tmp(39) := "0100" & "011" & "000000001010";
        tmp(40) := "0111" & "011" & "000000000000";
        tmp(41) := "1000" & "000" & "000000110001";
        tmp(42) := "0100" & "100" & "000000001011";
        tmp(43) := "0111" & "100" & "000000000000";
        tmp(44) := "1000" & "000" & "000000110101";
        tmp(45) := "0100" & "101" & "000000001100";
        tmp(46) := "0111" & "101" & "000000000000";
        tmp(47) := "1000" & "000" & "000000111001";
        tmp(48) := "1010" & "000" & "000000000111";
        tmp(49) := "0001" & "000" & "000000000001";
        tmp(50) := "0111" & "000" & "000000111100";
        tmp(51) := "1000" & "000" & "000000111101";
        tmp(52) := "1010" & "000" & "000000000111";
        tmp(53) := "0001" & "001" & "000000000001";
        tmp(54) := "0111" & "001" & "000000111100";
        tmp(55) := "1000" & "000" & "000000111111";
        tmp(56) := "1010" & "000" & "000000000111";
        tmp(57) := "0001" & "010" & "000000000001";
        tmp(58) := "0111" & "010" & "000000011000";
        tmp(59) := "1000" & "000" & "000001000001";
        tmp(60) := "1010" & "000" & "000000000111";
        tmp(61) := "0110" & "000" & "000000000000";
        tmp(62) := "1010" & "000" & "000000000111";
        tmp(63) := "0110" & "001" & "000000000000";
        tmp(64) := "1010" & "000" & "000000000111";
        tmp(65) := "0110" & "010" & "000000000000";
        tmp(66) := "1010" & "000" & "000000000111";

        RETURN tmp;
    END initMemory;

    SIGNAL memROM : blocoMemoria := initMemory;
BEGIN
    Dado <= memROM (to_integer(unsigned(Endereco)));
END ARCHITECTURE;